////////////////////////////////////////////////////////////////////////////////
// ECE 485/585: Microprocessor System Design
// Portland State University - Fall 2012 
// Final Project: 
// 
// File:		L_NEXT.v (Next Level Cache/Memory stub)
// Authors: 
// Description:
//
//
//
////////////////////////////////////////////////////////////////////////////////
module L_NEXT(
	// INPUTS
	input [25:0]  i_add_in,		// instruction cache address in
	input [25:0]  d_add_in		   // data cache address in
   );
	
endmodule
