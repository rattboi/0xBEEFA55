////////////////////////////////////////////////////////////////////////////////
// ECE 485/585: Microprocessor System Design
// Portland State University - Fall 2012 
// Final Project: 
// 
// File:		STATS.v (Statistics Module aka It's a series of counters)
// Authors: 
// Description:
//
//
//
////////////////////////////////////////////////////////////////////////////////
module STATS(
	// INPUTS
	input clk,				// clock may not be needed in this module
    input [3:0] n,			// mux to determine reads/writes
	input i_hit,       		// 
    input i_miss,        	// 
	input d_hit,       		// 
    input d_miss        	// 	
	
	// OUTPUTS 
	// none, will probably just use $display()
    );


endmodule
